///////////////////////////////////////////////////////////////////////////////
//     Copyright (c) 2025 Siliscale Consulting, LLC
// 
//    Licensed under the Apache License, Version 2.0 (the "License");
//    you may not use this file except in compliance with the License.
//    You may obtain a copy of the License at
// 
//        http://www.apache.org/licenses/LICENSE-2.0
// 
//    Unless required by applicable law or agreed to in writing, software
//    distributed under the License is distributed on an "AS IS" BASIS,
//    WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
//    See the License for the specific language governing permissions and
//    limitations under the License.
///////////////////////////////////////////////////////////////////////////////
//           _____          
//          /\    \         
//         /::\    \        
//        /::::\    \       
//       /::::::\    \      
//      /:::/\:::\    \     
//     /:::/__\:::\    \            Vendor      : Siliscale
//     \:::\   \:::\    \           Version     : 2025.1
//   ___\:::\   \:::\    \          Description : SVLib - Carry Save Adder (compressor) 4 to 2
//  /\   \:::\   \:::\    \ 
// /::\   \:::\   \:::\____\
// \:::\   \:::\   \::/    /
//  \:::\   \:::\   \/____/ 
//   \:::\   \:::\    \     
//    \:::\   \:::\____\    
//     \:::\  /:::/    /    
//      \:::\/:::/    /     
//       \::::::/    /      
//        \::::/    /       
//         \::/    /        
//          \/____/         
///////////////////////////////////////////////////////////////////////////////

module csa_4_2 #(
    parameter integer WIDTH = 32
) (
    input logic [WIDTH-1:0] in0,
    input logic [WIDTH-1:0] in1,
    input logic [WIDTH-1:0] in2,
    input logic [WIDTH-1:0] in3,

    output logic [WIDTH:0] sum,
    output logic [WIDTH:0] carry
);

  assign sum = {1'b0, in0 ^ in1 ^ in2 ^ in3} ^ {in3, 1'b0};  // Propagate

  assign carry = ({1'b0, (in0 & in1)}) |  // Generate
      ({1'b0, (in0 & in2)}) |  // Generate
      ({1'b0, in0} & {in3, 1'b0}) |  // Generate
      ({1'b0, in1} & {in3, 1'b0}) |  // Generate
      ({1'b0, in2} & {in3, 1'b0}) |  // Generate
      ({1'b0, in1 & in2});  // Generate





endmodule
